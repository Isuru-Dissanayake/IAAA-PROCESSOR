//module pc(
//
//input clock,
//output pc_out)
//
//
//
//end module
