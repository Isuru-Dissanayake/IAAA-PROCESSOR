module myInverter(
	input a,
	output out
	);
	
	assign out = -a;
	
endmodule