//
//
//
//
//module AC(           // ACCUMULATOR
//input clock,
//input [15:0] ALUOut,
//output [15:0] AC_out) 
//
//
//always @(posedge clock)
//begin
//
//end
//
//
//
//endmodule
